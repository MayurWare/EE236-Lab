Mayur Ware | 19D070070
*EE236 | Endsem | Q2 (a)
*NMOS Mobility
*Including NMOS model file
.include NMOSFET.txt

*Netlist
M1 D G GND GND NMOSFET L=0.4u W=1.2u AS={2*1.2u*0.4u} PS={2*1.2u+4*0.4u} AD={2*1.2u*0.4u} PD={2*1.2u+4*0.4u}    ;Definining NMOS 
V1 D1 D dc 0
Vd D1 GND dc 0.3
Vg G GND dc 0

*DC Analysis
.dc Vg 0.3 3.3 0.1
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot I(V1) vs V(G) ;ID vs VGS plot
.endc
.end
