Mayur Ware | 19D070070
*EE236 | Lab 6
*Id-Vgs Characteristics of NMOS
.include ALD1105N.txt               ;Including NMOS model file

*Netlist
M1 D G GND GND ALD1105N            ;Defining the NMOS Model Drain, Gate, Source, Body
*Vd D GND dc 200m
Vd D GND dc 5
Vg G GND dc 0

*DC Analysis
.dc Vg 0 5 0.01 
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2 
plot -I(Vd) vs V(G)             ;Id vs Vgs plot
plot sqrt(-I(Vd)) vs V(G)       ;sqrt(Id) vs Vgs plot
.endc
.end
