Mayur Ware | 19D070070
*EE236 | Midsem
*Voltage Regulator using Zener Diode
*Including BJT, Zener and Opamp model files
.include BZT52C18S.txt
.include bc547.txt
.include ua741.txt
*---------------------------------------

*-----------------------------------------
Vin 2 0 dc 21
Vsin 2 0 sin(0 18 50 0 0)
Rs 2 a 250k
Q1 2 c Out bc547a
X1 a b 2 0 c ua741
R1 Out b 16
R2 b 0 7k
X2 0 a DI_BZT52C18S

*Transient Analysis
.tran 10u 100m
*Control Commands
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot V(Out) vs V(2)
.endc
.end
