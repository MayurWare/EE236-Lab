Mayur Ware | 19D070070
*EE236 | Endsem | Q1 (a)
*Temperature Dependence of BJT
*Including BJT model file
.include bc547a.txt

*Netlist 
Q1 C B GND bc547a     ;Definining BJT 
V1 C2 C1 dc 0
V2 C2 GND dc 5
V3 B1 B dc 1
R2 B1 B 3k
R1 C C1 100

*DC Analysis
.dc V2 0 3 0.1 temp 25 55 10
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot I(V1) vs V(C)   ;Ic vs Vce plot
.endc
.end
