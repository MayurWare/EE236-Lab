Mayur Ware | 19D070070
*EE236 | Lab 2
*Voltage Regulator using Zener Diode
*Including BJT, Zener and Opamp model files
.include zener.txt
.include bc547.txt
.include ua741.txt
*---------------------------------------
*Bridge Rectifier using BAT85 Schottky Diode
*Including BAT85 Schottky Diode model file
.include schottky_BAT960.txt
*Bridge Rectifier
X1 1 2 BAT960
X2 0 1 BAT960
X3 3 2 BAT960
X4 0 3 BAT960
*Input Voltages
Vin 1 3 sin(0 16 50 0 0)
RL 2 0 1k
*Capacitor 
C1 2 0 1000u
*-----------------------------------------
Rs 2 a 52.64
Q1 2 c Out bc547a
X1 a b 2 0 c ua741
R1 Out b 6k
R2 b 0 10k
X2 0 a DI_1N4734A 

*Transient Analysis
.tran 10u 100m
*Control Commands
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot V(Out), V(2), V(3,1)
plot V(Out) vs V(3,1)
.endc
.end
