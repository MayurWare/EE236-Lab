Mayur Ware | 19D070070
*EE236 | Lab 5 | Part 1
*I-V Characteristics of PMOS
.include pmos.txt               ;Including PMOS model file

*Netlist
M1 D G GND GND ALD1107          ;Defining the PMOS Model Drain, Gate, Source, Body
Vd D GND dc 0
*Vg G GND dc -4
*Vg G GND dc -3.5
*Vg G GND dc -3
Vg G GND dc -2.5

*DC Analysis
.dc Vd -5 0 0.1 
.control
run
set color0 = white
set color1 = black
*set color2 = red 
*set color2 = blue
*set color2 = yellow
set color2 = green
set xbrushwidth = 2 
plot I(Vd) vs V(D)             ;Id vs Vds plot
plot abs((V(D))/(I(Vd)))        ;R_DS plot
.endc
.end
