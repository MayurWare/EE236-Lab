Mayur Ware | 19D070070
*EE236 | Midsem
*RN142S Analysis
*Including PIN Diode model file
.include Diode_1N914.txt
*Resistors 
R1 In 1 100
R2 1 0 1k
R3 3 0 100
*Diode 
D1 2 3 1N914
*Battery
Vin In 0 PULSE(0 5 0 0 0 0.5us 1us)
Vrd 1 2 dc 0
*Transient Analysis
.tran 1n 6u

.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
*Id vs Vd plot
let V = V(2) - V(3)
plot I(Vrd)
.endc
.end
