Mayur Ware | 19D070070
*EE236 | Midsem
*Temperature Dependence of Zener Diode
*Including Zener Diode Model File
.include BZT52C18S.txt
*Resistors 
R1 In 1 100
R2 1 0 1k
R3 3 0 100
*Diode 
X1 3 2 DI_BZT52C18S
*Battery
Vin In 0 dc 0.01
Vbl 1 2 dc 0
*DC Analysis
.dc vin 0 19.31 19.31 temp 20 80 10

.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
*Id vs Vd plot
let V = V(2) - V(3)
plot V
.endc
.end
