Mayur Ware | 19D070070
*EE236 | Lab 0 | Exercise 2
*Bridge Rectifier analysis
*Including Diode model file
.include Diode_1N914.txt
*Bridge Rectifier
D1 1 2 1N914
D2 0 1 1N914
D3 3 2 1N914
D4 0 3 1N914
*Load Resistor
R1 2 0 1k
*Input Voltages
Vin 1 3 sin(0 12 50 0 0)
*Transient Analysis
.tran 10u 100m
*Control Commands
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
let V_input = V(1) - V(3)
plot V(2) V_input
plot V(2) vs V_input
.endc
.end