Mayur Ware | 19D070070
*EE236 | Quiz 1 | Q3
*Including Model files
.include schottky_bat85.cir
.include TL071.cir

*Netlist
R1 1 3 10k
R2 2 3 1k
Rf 3 4 1k
Rfb 5 Out 150k
Cfb 5 Out 100p
X1 0 3 a b 4 TL071
X2 0 5 c d Out TL071
X3 5 4 BAT85

*Voltages 
Vdc GND 2 dc 0.01
Vsin 0 1 sin(0 1 100k 0 0)
Va GND1 a dc 15
Vb b GND2 dc 15
Vc GND3 c dc 15
Vd d GND4 dc 15

*DC Analysis
.dc Vdc 0 5 0.01
*Control Commands
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2
plot V(4)
plot V(Out) vs V(4)
.endc
.end
