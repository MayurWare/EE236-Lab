Mayur Ware | 19D070070
*EE236 | Lab 3
*Including Model files
.include TL071.cir
.include Solar_Cell.cir

*Netlist
R1 1 3 10k
R2 2 3 1k
Rf 3 4 1k
Rfb 5 Out 150k
Cfb 5 Out 100p
X1 0 3 a b 4 TL071
X2 0 5 c d Out TL071
X3 5 4 solar_cell IL_val = 0e-3

*Voltages 
Vdc GND 2 dc 0.01
Vsin 0 1 sin(0 1 100k 0 0)
Va GND a dc 15
Vb GND b dc -15
Vc GND c dc 15
Vd GND d dc -15

*DC Analysis
.dc Vdc 0 2 0.01
*Control Commands
.control
run
set color0 = white
set color1 = black
set color2 = blue
set color3 = red
set xbrushwidth = 2

let C=4.7e-9
let R=10k
let w=6.28k
let Cdut = (V(Out)*C*sqrt(1+1/(w*C*R)^2)/V(4,5)
.endc
.end
